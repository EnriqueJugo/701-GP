-- megafunction wizard: %LPM_MUX%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: LPM_MUX 

-- ============================================================
-- File Name: mux_2.vhd
-- Megafunction Name(s):
-- 			LPM_MUX
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 18.1.0 Build 625 09/12/2018 SJ Standard Edition
-- ************************************************************


--Copyright (C) 2018  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel FPGA IP License Agreement, or other applicable license
--agreement, including, without limitation, that your use is for
--the sole purpose of programming logic devices manufactured by
--Intel and sold by Intel or its authorized distributors.  Please
--refer to the applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY lpm;
USE lpm.lpm_components.all;

ENTITY mux_2 IS
	PORT
	(
		data0x		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		data1x		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		data2x		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		data3x		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		sel		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
	);
END mux_2;


ARCHITECTURE SYN OF mux_2 IS

--	type STD_LOGIC_2D is array (NATURAL RANGE <>, NATURAL RANGE <>) of STD_LOGIC;

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_2D (3 DOWNTO 0, 15 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (15 DOWNTO 0);

BEGIN
	sub_wire4    <= data0x(15 DOWNTO 0);
	sub_wire3    <= data1x(15 DOWNTO 0);
	sub_wire2    <= data2x(15 DOWNTO 0);
	sub_wire0    <= data3x(15 DOWNTO 0);
	sub_wire1(3, 0)    <= sub_wire0(0);
	sub_wire1(3, 1)    <= sub_wire0(1);
	sub_wire1(3, 2)    <= sub_wire0(2);
	sub_wire1(3, 3)    <= sub_wire0(3);
	sub_wire1(3, 4)    <= sub_wire0(4);
	sub_wire1(3, 5)    <= sub_wire0(5);
	sub_wire1(3, 6)    <= sub_wire0(6);
	sub_wire1(3, 7)    <= sub_wire0(7);
	sub_wire1(3, 8)    <= sub_wire0(8);
	sub_wire1(3, 9)    <= sub_wire0(9);
	sub_wire1(3, 10)    <= sub_wire0(10);
	sub_wire1(3, 11)    <= sub_wire0(11);
	sub_wire1(3, 12)    <= sub_wire0(12);
	sub_wire1(3, 13)    <= sub_wire0(13);
	sub_wire1(3, 14)    <= sub_wire0(14);
	sub_wire1(3, 15)    <= sub_wire0(15);
	sub_wire1(2, 0)    <= sub_wire2(0);
	sub_wire1(2, 1)    <= sub_wire2(1);
	sub_wire1(2, 2)    <= sub_wire2(2);
	sub_wire1(2, 3)    <= sub_wire2(3);
	sub_wire1(2, 4)    <= sub_wire2(4);
	sub_wire1(2, 5)    <= sub_wire2(5);
	sub_wire1(2, 6)    <= sub_wire2(6);
	sub_wire1(2, 7)    <= sub_wire2(7);
	sub_wire1(2, 8)    <= sub_wire2(8);
	sub_wire1(2, 9)    <= sub_wire2(9);
	sub_wire1(2, 10)    <= sub_wire2(10);
	sub_wire1(2, 11)    <= sub_wire2(11);
	sub_wire1(2, 12)    <= sub_wire2(12);
	sub_wire1(2, 13)    <= sub_wire2(13);
	sub_wire1(2, 14)    <= sub_wire2(14);
	sub_wire1(2, 15)    <= sub_wire2(15);
	sub_wire1(1, 0)    <= sub_wire3(0);
	sub_wire1(1, 1)    <= sub_wire3(1);
	sub_wire1(1, 2)    <= sub_wire3(2);
	sub_wire1(1, 3)    <= sub_wire3(3);
	sub_wire1(1, 4)    <= sub_wire3(4);
	sub_wire1(1, 5)    <= sub_wire3(5);
	sub_wire1(1, 6)    <= sub_wire3(6);
	sub_wire1(1, 7)    <= sub_wire3(7);
	sub_wire1(1, 8)    <= sub_wire3(8);
	sub_wire1(1, 9)    <= sub_wire3(9);
	sub_wire1(1, 10)    <= sub_wire3(10);
	sub_wire1(1, 11)    <= sub_wire3(11);
	sub_wire1(1, 12)    <= sub_wire3(12);
	sub_wire1(1, 13)    <= sub_wire3(13);
	sub_wire1(1, 14)    <= sub_wire3(14);
	sub_wire1(1, 15)    <= sub_wire3(15);
	sub_wire1(0, 0)    <= sub_wire4(0);
	sub_wire1(0, 1)    <= sub_wire4(1);
	sub_wire1(0, 2)    <= sub_wire4(2);
	sub_wire1(0, 3)    <= sub_wire4(3);
	sub_wire1(0, 4)    <= sub_wire4(4);
	sub_wire1(0, 5)    <= sub_wire4(5);
	sub_wire1(0, 6)    <= sub_wire4(6);
	sub_wire1(0, 7)    <= sub_wire4(7);
	sub_wire1(0, 8)    <= sub_wire4(8);
	sub_wire1(0, 9)    <= sub_wire4(9);
	sub_wire1(0, 10)    <= sub_wire4(10);
	sub_wire1(0, 11)    <= sub_wire4(11);
	sub_wire1(0, 12)    <= sub_wire4(12);
	sub_wire1(0, 13)    <= sub_wire4(13);
	sub_wire1(0, 14)    <= sub_wire4(14);
	sub_wire1(0, 15)    <= sub_wire4(15);
	result    <= sub_wire5(15 DOWNTO 0);

	LPM_MUX_component : LPM_MUX
	GENERIC MAP (
		lpm_size => 4,
		lpm_type => "LPM_MUX",
		lpm_width => 16,
		lpm_widths => 2
	)
	PORT MAP (
		data => sub_wire1,
		sel => sel,
		result => sub_wire5
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: new_diagram STRING "1"
-- Retrieval info: LIBRARY: lpm lpm.lpm_components.all
-- Retrieval info: CONSTANT: LPM_SIZE NUMERIC "4"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MUX"
-- Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "16"
-- Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "2"
-- Retrieval info: USED_PORT: data0x 0 0 16 0 INPUT NODEFVAL "data0x[15..0]"
-- Retrieval info: USED_PORT: data1x 0 0 16 0 INPUT NODEFVAL "data1x[15..0]"
-- Retrieval info: USED_PORT: data2x 0 0 16 0 INPUT NODEFVAL "data2x[15..0]"
-- Retrieval info: USED_PORT: data3x 0 0 16 0 INPUT NODEFVAL "data3x[15..0]"
-- Retrieval info: USED_PORT: result 0 0 16 0 OUTPUT NODEFVAL "result[15..0]"
-- Retrieval info: USED_PORT: sel 0 0 2 0 INPUT NODEFVAL "sel[1..0]"
-- Retrieval info: CONNECT: @data 1 0 16 0 data0x 0 0 16 0
-- Retrieval info: CONNECT: @data 1 1 16 0 data1x 0 0 16 0
-- Retrieval info: CONNECT: @data 1 2 16 0 data2x 0 0 16 0
-- Retrieval info: CONNECT: @data 1 3 16 0 data3x 0 0 16 0
-- Retrieval info: CONNECT: @sel 0 0 2 0 sel 0 0 2 0
-- Retrieval info: CONNECT: result 0 0 16 0 @result 0 0 16 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux_2.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux_2.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux_2.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux_2.bsf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux_2_inst.vhd FALSE
-- Retrieval info: LIB_FILE: lpm
